CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 2850 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
76 E:\2.2 - Study materials\CSE 210 (Digital Logic & System Design LAB)\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
56
13 Logic Switch~
5 376 3202 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44592 0
0
13 Logic Switch~
5 357 3103 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44592 0
0
13 Logic Switch~
5 213 3056 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44592 0
0
13 Logic Switch~
5 256 2865 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.90018e-315 0
0
13 Logic Switch~
5 253 2921 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
0 -25 7 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90018e-315 0
0
13 Logic Switch~
5 165 2042 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-7 -21 7 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.90018e-315 0
0
13 Logic Switch~
5 57 2036 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-2 -19 12 -11
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.90018e-315 0
0
13 Logic Switch~
5 112 2039 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90018e-315 0
0
13 Logic Switch~
5 136 1449 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
44592 0
0
13 Logic Switch~
5 130 1376 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
44592 1
0
13 Logic Switch~
5 127 1294 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
44592 2
0
13 Logic Switch~
5 273 1006 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.90018e-315 0
0
13 Logic Switch~
5 235 902 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
5.90018e-315 5.26354e-315
0
13 Logic Switch~
5 167 878 0 1 11
0 40
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.90018e-315 5.30499e-315
0
13 Logic Switch~
5 87 111 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -18 8 -10
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3835 0 0
2
5.90018e-315 5.32571e-315
0
13 Logic Switch~
5 95 50 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3670 0 0
2
5.90018e-315 5.34643e-315
0
13 Logic Switch~
5 216 412 0 1 11
0 44
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 Cin
-9 -30 12 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.90018e-315 5.3568e-315
0
13 Logic Switch~
5 173 410 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9323 0 0
2
5.90018e-315 5.36716e-315
0
13 Logic Switch~
5 131 410 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
317 0 0
2
5.90018e-315 5.37752e-315
0
9 2-In AND~
219 398 2358 0 3 22
0 7 6 11
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3108 0 0
2
44592.1 0
0
9 2-In AND~
219 321 2486 0 3 22
0 3 5 25
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
4299 0 0
2
44592.1 0
0
9 2-In AND~
219 267 2233 0 3 22
0 3 4 2
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
9672 0 0
2
44592.1 0
0
9 2-In AND~
219 665 2133 0 3 22
0 13 12 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
7876 0 0
2
44592.1 0
0
8 2-In OR~
219 885 2246 0 3 22
0 9 10 8
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
6369 0 0
2
44592 0
0
8 2-In OR~
219 587 2517 0 3 22
0 25 5 10
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
9172 0 0
2
44592 0
0
8 2-In OR~
219 508 2234 0 3 22
0 2 11 12
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
7100 0 0
2
44592 0
0
8 2-In OR~
219 320 2090 0 3 22
0 14 5 13
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3820 0 0
2
44592 0
0
8 2-In OR~
219 426 2898 0 3 22
0 17 16 15
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
1 -25 15 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
7678 0 0
2
44592 0
0
9 2-In AND~
219 542 3171 0 3 22
0 21 22 18
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
961 0 0
2
44592 0
0
9 2-In AND~
219 495 3082 0 3 22
0 23 24 19
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3178 0 0
2
44592 0
0
8 2-In OR~
219 649 3073 0 3 22
0 19 18 20
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
1 -25 15 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3409 0 0
2
44592 0
0
9 Inverter~
13 288 3168 0 2 22
0 23 21
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
3951 0 0
2
44592 0
0
14 Logic Display~
6 781 3066 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
44592 0
0
14 Logic Display~
6 542 2867 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.90018e-315 0
0
14 Logic Display~
6 1014 2170 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
5.90018e-315 0
0
9 Inverter~
13 258 2398 0 2 22
0 4 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9442 0 0
2
5.90018e-315 0
0
14 Logic Display~
6 833 1337 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
44592 3
0
8 2-In OR~
219 767 1372 0 3 22
0 28 27 26
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9968 0 0
2
44592 4
0
8 2-In OR~
219 669 1280 0 3 22
0 30 29 28
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9281 0 0
2
44592 5
0
9 2-In AND~
219 354 1456 0 3 22
0 31 32 27
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
8464 0 0
2
44592 6
0
9 2-In AND~
219 338 1357 0 3 22
0 33 32 29
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7168 0 0
2
44592 7
0
9 2-In AND~
219 338 1277 0 3 22
0 31 33 30
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3171 0 0
2
44592 8
0
8 2-In OR~
219 610 932 0 3 22
0 37 35 34
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OD
1 -25 15 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
4139 0 0
2
5.90018e-315 5.38788e-315
0
9 2-In AND~
219 420 1107 0 3 22
0 39 38 35
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
6435 0 0
2
5.90018e-315 5.39306e-315
0
9 2-In AND~
219 454 884 0 3 22
0 40 36 37
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 ANC
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5283 0 0
2
5.90018e-315 5.39824e-315
0
9 Inverter~
13 222 960 0 2 22
0 40 39
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
6874 0 0
2
5.90018e-315 5.40342e-315
0
14 Logic Display~
6 921 840 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.90018e-315 5.4086e-315
0
14 Logic Display~
6 1082 517 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.90018e-315 5.41378e-315
0
8 2-In OR~
219 754 661 0 3 22
0 43 42 41
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
969 0 0
2
5.90018e-315 5.41896e-315
0
9 2-In AND~
219 642 702 0 3 22
0 45 44 42
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8402 0 0
2
5.90018e-315 5.42414e-315
0
14 Logic Display~
6 696 394 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -20 7 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.90018e-315 5.42933e-315
0
9 2-In XOR~
219 560 447 0 3 22
0 45 44 48
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4292 0 0
2
5.90018e-315 5.43192e-315
0
9 2-In XOR~
219 360 395 0 3 22
0 47 46 45
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6118 0 0
2
5.90018e-315 5.43451e-315
0
14 Logic Display~
6 1115 196 0 1 2
10 49
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.90018e-315 5.4371e-315
0
8 2-In OR~
219 862 164 0 3 22
0 51 50 49
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OC
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6357 0 0
2
5.90018e-315 5.43969e-315
0
9 2-In AND~
219 630 540 0 3 22
0 47 46 43
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
319 0 0
2
5.90018e-315 5.44228e-315
0
63
1 3 2 0 0 4224 0 26 22 0 0 4
495 2225
296 2225
296 2233
288 2233
1 0 3 0 0 4096 0 22 0 0 4 2
243 2224
57 2224
2 0 4 0 0 4096 0 22 0 0 27 2
243 2242
165 2242
1 1 3 0 0 8320 0 21 7 0 0 3
297 2477
57 2477
57 2048
2 0 5 0 0 4096 0 21 0 0 29 2
297 2495
112 2495
2 2 6 0 0 4224 0 20 36 0 0 4
374 2367
287 2367
287 2398
279 2398
1 0 7 0 0 4224 0 20 0 0 0 2
374 2349
57 2349
1 3 8 0 0 8320 0 35 24 0 0 3
1014 2188
1014 2246
918 2246
1 3 9 0 0 4224 0 24 23 0 0 4
872 2237
694 2237
694 2133
686 2133
2 3 10 0 0 8320 0 24 25 0 0 4
872 2255
628 2255
628 2517
620 2517
2 3 11 0 0 8320 0 26 20 0 0 4
495 2243
427 2243
427 2358
419 2358
2 3 12 0 0 4224 0 23 26 0 0 4
641 2142
549 2142
549 2234
541 2234
1 3 13 0 0 4224 0 23 27 0 0 4
641 2124
361 2124
361 2090
353 2090
2 0 5 0 0 4096 0 27 0 0 29 2
307 2099
112 2099
1 0 14 0 0 4224 0 27 0 0 0 2
307 2081
57 2081
1 3 15 0 0 8320 0 34 28 0 0 3
542 2885
542 2898
459 2898
2 1 16 0 0 4224 0 28 5 0 0 4
413 2907
274 2907
274 2921
265 2921
1 1 17 0 0 4224 0 28 4 0 0 4
413 2889
277 2889
277 2865
268 2865
2 3 18 0 0 8320 0 31 29 0 0 4
636 3082
571 3082
571 3171
563 3171
1 3 19 0 0 4224 0 31 30 0 0 4
636 3064
524 3064
524 3082
516 3082
3 1 20 0 0 4224 0 31 33 0 0 5
682 3073
769 3073
769 3092
781 3092
781 3084
1 2 21 0 0 4224 0 29 32 0 0 4
518 3162
317 3162
317 3168
309 3168
2 1 22 0 0 4224 0 29 1 0 0 4
518 3180
397 3180
397 3202
388 3202
1 0 23 0 0 8192 0 32 0 0 26 3
273 3168
267 3168
267 3073
2 1 24 0 0 4224 0 30 2 0 0 4
471 3091
378 3091
378 3103
369 3103
1 1 23 0 0 4224 0 30 3 0 0 4
471 3073
234 3073
234 3056
225 3056
1 1 4 0 0 8320 0 36 6 0 0 3
243 2398
165 2398
165 2054
1 3 25 0 0 8320 0 25 21 0 0 6
574 2508
574 2510
350 2510
350 2489
342 2489
342 2486
2 1 5 0 0 12416 0 25 8 0 0 4
574 2526
574 2528
112 2528
112 2051
3 1 26 0 0 4224 0 38 37 0 0 3
800 1372
833 1372
833 1355
2 3 27 0 0 4224 0 38 40 0 0 4
754 1381
383 1381
383 1456
375 1456
3 1 28 0 0 20608 0 39 38 0 0 6
702 1280
723 1280
723 1338
665 1338
665 1363
754 1363
3 2 29 0 0 4224 0 41 39 0 0 4
359 1357
648 1357
648 1289
656 1289
3 1 30 0 0 4224 0 42 39 0 0 4
359 1277
648 1277
648 1271
656 1271
0 1 31 0 0 4096 0 0 40 40 0 3
267 1294
267 1447
330 1447
0 2 32 0 0 4096 0 0 41 38 0 3
238 1449
238 1366
314 1366
0 2 33 0 0 4096 0 0 42 39 0 3
241 1376
241 1286
314 1286
1 2 32 0 0 4224 0 9 40 0 0 4
148 1449
322 1449
322 1465
330 1465
1 1 33 0 0 4224 0 10 41 0 0 4
142 1376
306 1376
306 1348
314 1348
1 1 31 0 0 4224 0 11 42 0 0 4
139 1294
306 1294
306 1268
314 1268
3 1 34 0 0 12416 0 43 47 0 0 5
643 932
639 932
639 917
921 917
921 858
2 3 35 0 0 8320 0 43 44 0 0 4
597 941
447 941
447 1107
441 1107
1 2 36 0 0 4224 0 13 45 0 0 4
247 902
341 902
341 893
430 893
3 1 37 0 0 12416 0 45 43 0 0 4
475 884
516 884
516 923
597 923
2 1 38 0 0 8320 0 44 12 0 0 4
396 1116
294 1116
294 1006
285 1006
2 1 39 0 0 8320 0 46 44 0 0 4
243 960
363 960
363 1098
396 1098
0 1 40 0 0 4096 0 0 46 48 0 3
209 878
209 960
207 960
1 1 40 0 0 4224 0 14 45 0 0 4
179 878
341 878
341 875
430 875
1 3 41 0 0 4224 0 48 49 0 0 3
1082 535
787 535
787 661
3 2 42 0 0 12416 0 50 49 0 0 4
663 702
679 702
679 670
741 670
3 1 43 0 0 8320 0 56 49 0 0 4
651 540
679 540
679 652
741 652
0 2 44 0 0 8192 0 0 50 57 0 3
379 510
379 711
618 711
0 1 45 0 0 8320 0 0 50 58 0 3
413 493
413 693
618 693
2 1 46 0 0 4224 0 56 18 0 0 3
606 549
173 549
173 422
1 1 47 0 0 4224 0 56 19 0 0 3
606 531
131 531
131 422
1 3 48 0 0 8320 0 51 52 0 0 3
696 412
696 447
593 447
1 2 44 0 0 12416 0 17 52 0 0 5
216 424
217 424
217 510
544 510
544 456
1 3 45 0 0 0 0 52 53 0 0 6
544 438
413 438
413 493
395 493
395 395
393 395
2 0 46 0 0 0 0 53 0 0 54 5
344 404
344 426
188 426
188 477
173 477
1 0 47 0 0 0 0 53 0 0 55 5
344 386
344 373
146 373
146 459
131 459
3 1 49 0 0 8320 0 55 54 0 0 3
895 164
895 214
1115 214
1 2 50 0 0 8320 0 15 55 0 0 5
99 111
99 291
749 291
749 173
849 173
1 1 51 0 0 8320 0 16 55 0 0 5
107 50
107 48
750 48
750 155
849 155
67
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
239 2096 300 2120
249 2104 289 2120
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
475 2524 536 2548
485 2532 525 2548
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
474 2483 535 2507
484 2491 524 2507
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
625 2463 686 2487
635 2471 675 2487
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
336 2459 397 2483
346 2467 386 2483
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
238 2493 299 2517
248 2501 288 2517
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
236 2452 297 2476
246 2460 286 2476
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
253 2394 314 2418
263 2402 303 2418
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
190 2396 251 2420
200 2404 240 2420
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
422 2330 483 2354
432 2338 472 2354
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
327 2364 388 2388
337 2372 377 2388
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
327 2322 388 2346
337 2330 377 2346
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
544 2214 605 2238
554 2222 594 2238
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
437 2238 498 2262
447 2246 487 2262
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
444 2199 505 2223
454 2207 494 2223
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
190 2238 251 2262
200 2246 240 2262
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
187 2199 248 2223
197 2207 237 2223
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
301 2199 362 2223
311 2207 351 2223
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
929 2217 990 2241
939 2225 979 2241
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
795 2253 856 2277
805 2261 845 2277
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
797 2207 858 2231
807 2215 847 2231
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
677 2107 738 2131
687 2115 727 2131
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
584 2136 645 2160
594 2144 634 2160
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
584 2094 645 2118
594 2102 634 2118
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
338 2062 399 2086
348 2070 388 2086
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
239 2054 300 2078
249 2062 289 2078
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
660 1856 761 1880
670 1864 750 1880
10 B I BEFORE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
819 251 864 275
829 259 853 275
3 A+C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
33 22 58 46
41 30 49 46
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
73 772 102 796
83 780 91 796
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
701 363 746 387
711 371 735 387
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1097 483 1158 507
1107 491 1147 507
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
924 533 985 557
934 541 974 557
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
685 620 746 644
695 628 735 644
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
690 665 743 689
700 673 732 689
4 pin2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
651 514 712 538
661 522 701 538
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
650 699 711 723
660 707 700 723
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
553 668 614 692
563 676 603 692
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
535 507 596 531
545 515 585 531
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
535 542 596 566
545 550 585 566
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
552 704 613 728
562 712 602 728
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
620 417 681 441
630 425 670 441
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
463 485 524 509
473 493 513 509
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
458 412 519 436
468 420 508 436
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
380 368 441 392
390 376 430 392
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
235 349 296 373
245 357 285 373
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
240 423 301 447
250 431 290 447
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
429 2927 490 2951
439 2935 479 2951
5 Y=A+C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
487 1438 580 1462
497 1446 569 1462
9  AB+BC+AC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
472 2873 533 2897
482 2881 522 2897
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
318 2861 379 2885
328 2869 368 2885
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
320 2901 381 2925
330 2909 370 2925
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
767 1317 828 1341
777 1325 817 1341
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
690 1338 751 1362
700 1346 740 1362
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
699 1378 760 1402
709 1386 749 1402
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
694 1252 755 1276
704 1260 744 1276
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
574 1254 635 1278
584 1262 624 1278
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
577 1332 638 1356
587 1340 627 1356
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
360 1250 421 1274
370 1258 410 1274
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
368 1331 429 1355
378 1339 418 1355
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
362 1456 423 1480
372 1464 412 1480
5 pin 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
240 1447 301 1471
250 1455 290 1471
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
268 1419 329 1443
278 1427 318 1443
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
266 1372 327 1396
276 1380 316 1396
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
179 1347 240 1371
189 1355 229 1371
5 pin 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
292 1290 353 1314
302 1298 342 1314
5 pin 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
174 1265 235 1289
184 1273 224 1289
5 pin 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
