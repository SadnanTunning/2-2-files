CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 587 193 0 1 11
0 2
0
0 0 21360 0
2 0V
-32 -5 -18 3
1 R
24 -12 31 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44609.9 0
0
13 Logic Switch~
5 586 101 0 1 11
0 3
0
0 0 21360 0
2 0V
-32 0 -18 8
1 S
26 -10 33 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44609.9 1
0
13 Logic Switch~
5 113 174 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -7 -16 1
1 R
21 -11 28 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44609.9 2
0
13 Logic Switch~
5 111 96 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-33 -2 -19 6
1 S
23 -14 30 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44609.9 3
0
14 Logic Display~
6 814 168 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
44609.9 4
0
14 Logic Display~
6 813 94 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44609.9 5
0
14 Logic Display~
6 372 146 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
44609.9 6
0
14 Logic Display~
6 372 88 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
44609.9 7
0
10 2-In NAND~
219 247 105 0 3 22
0 7 5 4
0
0 0 624 0
4 7400
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
5.9002e-315 0
0
10 2-In NAND~
219 247 165 0 3 22
0 4 6 5
0
0 0 624 0
4 7400
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
5.9002e-315 5.26354e-315
0
9 2-In NOR~
219 702 111 0 3 22
0 3 9 8
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 NOR
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3472 0 0
2
5.9002e-315 5.30499e-315
0
9 2-In NOR~
219 704 185 0 3 22
0 8 2 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 NOR
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9998 0 0
2
5.9002e-315 5.32571e-315
0
12
1 2 2 0 0 8320 0 1 12 0 0 3
599 193
599 194
691 194
1 1 3 0 0 8320 0 2 11 0 0 3
598 101
598 102
689 102
0 1 4 0 0 8320 0 0 10 6 0 5
305 105
305 128
159 128
159 156
223 156
2 0 5 0 0 12416 0 9 0 0 5 5
223 114
174 114
174 138
305 138
305 165
3 1 5 0 0 0 0 10 7 0 0 3
274 165
372 165
372 164
3 1 4 0 0 0 0 9 8 0 0 4
274 105
305 105
305 106
372 106
1 2 6 0 0 4224 0 3 10 0 0 2
125 174
223 174
1 1 7 0 0 4224 0 4 9 0 0 2
123 96
223 96
1 0 8 0 0 12416 0 12 0 0 12 5
691 176
646 176
646 141
764 141
764 111
2 0 9 0 0 12416 0 11 0 0 11 5
689 120
627 120
627 155
767 155
767 185
3 1 9 0 0 0 0 12 5 0 0 3
743 185
814 185
814 186
3 1 8 0 0 0 0 11 6 0 0 3
741 111
813 111
813 112
18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
665 192 690 213
673 199 681 214
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
663 155 690 176
672 162 680 177
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
763 186 790 207
772 193 780 208
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
664 115 691 136
673 121 681 136
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
663 75 690 96
672 82 680 97
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
768 87 795 108
777 93 785 108
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
321 146 346 167
329 153 337 168
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
186 168 211 189
194 175 202 190
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
185 134 210 155
193 141 201 156
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
317 79 344 100
326 86 334 101
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
186 93 211 114
194 99 202 114
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
186 72 213 93
195 78 203 93
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
828 75 865 99
838 83 854 99
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
381 124 418 148
391 132 407 148
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
838 162 867 186
848 170 856 186
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
832 89 861 113
842 97 850 113
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
385 140 414 164
395 148 403 164
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
381 80 410 104
391 88 399 104
1 Q
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
