CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
65
13 Logic Switch~
5 653 1157 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44599.9 0
0
13 Logic Switch~
5 652 1083 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44599.9 1
0
13 Logic Switch~
5 89 1188 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44599.9 2
0
13 Logic Switch~
5 90 1109 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44599.9 3
0
13 Logic Switch~
5 718 958 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90019e-315 0
0
13 Logic Switch~
5 711 915 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90019e-315 5.26354e-315
0
13 Logic Switch~
5 112 962 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90019e-315 5.30499e-315
0
13 Logic Switch~
5 111 923 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90019e-315 5.32571e-315
0
13 Logic Switch~
5 662 733 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90019e-315 5.34643e-315
0
13 Logic Switch~
5 667 670 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90019e-315 5.3568e-315
0
13 Logic Switch~
5 94 776 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -16 9 -8
3 V12
-5 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90019e-315 5.36716e-315
0
13 Logic Switch~
5 103 703 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90019e-315 5.37752e-315
0
13 Logic Switch~
5 675 345 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90019e-315 5.38788e-315
0
13 Logic Switch~
5 140 468 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.90019e-315 5.39306e-315
0
13 Logic Switch~
5 677 481 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.90019e-315 5.39824e-315
0
13 Logic Switch~
5 677 561 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.90019e-315 5.40342e-315
0
13 Logic Switch~
5 665 248 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -15 8 -7
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.90019e-315 5.4086e-315
0
13 Logic Switch~
5 703 125 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.90019e-315 5.41378e-315
0
13 Logic Switch~
5 138 575 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.90019e-315 5.41896e-315
0
13 Logic Switch~
5 166 327 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3108 0 0
2
5.90019e-315 5.42414e-315
0
13 Logic Switch~
5 162 273 0 10 11
0 52 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4299 0 0
2
5.90019e-315 5.42933e-315
0
13 Logic Switch~
5 158 123 0 10 11
0 53 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9672 0 0
2
5.90019e-315 5.43192e-315
0
5 4001~
219 797 931 0 3 22
0 10 9 5
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 10 0
1 U
7876 0 0
2
44599.9 4
0
5 4011~
219 209 936 0 3 22
0 8 7 6
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 7 0
1 U
6369 0 0
2
44599.9 5
0
5 4001~
219 952 1111 0 3 22
0 17 17 15
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 8 0
1 U
9172 0 0
2
44599.9 6
0
5 4001~
219 833 1115 0 3 22
0 20 19 17
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 8 0
1 U
7100 0 0
2
44599.9 7
0
5 4001~
219 732 1157 0 3 22
0 12 12 19
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 8 0
1 U
3820 0 0
2
44599.9 8
0
5 4001~
219 732 1088 0 3 22
0 11 11 20
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 8 0
1 U
7678 0 0
2
44599.9 9
0
5 4011~
219 356 1137 0 3 22
0 18 18 16
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 7 0
1 U
961 0 0
2
44599.9 10
0
5 4011~
219 254 1139 0 3 22
0 22 21 18
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 7 0
1 U
3178 0 0
2
44599.9 11
0
5 4011~
219 161 1115 0 3 22
0 14 14 22
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 7 0
1 U
3409 0 0
2
44599.9 12
0
5 4011~
219 172 1179 0 3 22
0 13 13 21
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 3 0
1 U
3951 0 0
2
44599.9 13
0
5 4001~
219 1045 681 0 3 22
0 24 24 23
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 6 0
1 U
8885 0 0
2
5.90019e-315 5.43451e-315
0
5 4001~
219 938 676 0 3 22
0 26 25 24
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 6 0
1 U
3780 0 0
2
5.90019e-315 5.4371e-315
0
5 4001~
219 849 715 0 3 22
0 4 3 25
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 6 0
1 U
9265 0 0
2
5.90019e-315 5.43969e-315
0
5 4001~
219 839 650 0 3 22
0 2 4 26
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 5 0
1 U
9442 0 0
2
5.90019e-315 5.44228e-315
0
5 4001~
219 734 699 0 3 22
0 2 3 4
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 5 0
1 U
9424 0 0
2
5.90019e-315 5.44487e-315
0
5 4001~
219 924 304 0 3 22
0 40 39 41
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 5 0
1 U
9968 0 0
2
5.90019e-315 5.44746e-315
0
5 4001~
219 922 513 0 3 22
0 35 35 36
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 5 0
1 U
9281 0 0
2
5.90019e-315 5.45005e-315
0
5 4001~
219 777 510 0 3 22
0 34 33 35
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 4 0
1 U
8464 0 0
2
5.90019e-315 5.45264e-315
0
5 4001~
219 754 341 0 3 22
0 38 38 39
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 4 0
1 U
7168 0 0
2
5.90019e-315 5.45523e-315
0
5 4001~
219 739 246 0 3 22
0 37 37 40
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 4 0
1 U
3171 0 0
2
5.90019e-315 5.45782e-315
0
5 4001~
219 826 118 0 3 22
0 42 42 43
0
0 0 624 0
4 4001
-14 -24 14 -16
3 NOR
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 4 0
1 U
4139 0 0
2
5.90019e-315 5.46041e-315
0
14 Logic Display~
6 1058 282 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
5.90019e-315 5.463e-315
0
14 Logic Display~
6 1020 87 0 1 2
10 43
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.90019e-315 5.46559e-315
0
14 Logic Display~
6 1121 660 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
5.90019e-315 5.46818e-315
0
14 Logic Display~
6 418 901 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.90019e-315 5.47077e-315
0
14 Logic Display~
6 1046 1095 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.90019e-315 5.47207e-315
0
14 Logic Display~
6 457 504 0 1 2
10 44
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.90019e-315 5.47336e-315
0
14 Logic Display~
6 489 715 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.90019e-315 5.47466e-315
0
14 Logic Display~
6 1017 483 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.90019e-315 5.47595e-315
0
14 Logic Display~
6 1017 903 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
5.90019e-315 5.47725e-315
0
14 Logic Display~
6 430 1102 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.90019e-315 5.47854e-315
0
14 Logic Display~
6 488 288 0 1 2
10 49
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.90019e-315 5.47984e-315
0
5 4011~
219 223 567 0 3 22
0 47 47 46
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 3 0
1 U
6357 0 0
2
5.90019e-315 5.48113e-315
0
5 4011~
219 347 529 0 3 22
0 45 46 44
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 3 0
1 U
319 0 0
2
5.90019e-315 5.48243e-315
0
5 4011~
219 267 776 0 3 22
0 32 31 28
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 2 0
1 U
3976 0 0
2
5.90019e-315 5.48372e-315
0
5 4011~
219 171 743 0 3 22
0 30 31 32
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 2 0
1 U
7634 0 0
2
5.90019e-315 5.48502e-315
0
5 4011~
219 368 745 0 3 22
0 29 28 27
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 2 0
1 U
523 0 0
2
5.90019e-315 5.48631e-315
0
5 4011~
219 266 706 0 3 22
0 30 32 29
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
6748 0 0
2
5.90019e-315 5.48761e-315
0
5 4011~
219 220 487 0 3 22
0 48 48 45
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 1 0
1 U
6901 0 0
2
5.90019e-315 5.4889e-315
0
5 4011~
219 377 293 0 3 22
0 50 50 49
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
842 0 0
2
5.90019e-315 5.4902e-315
0
5 4011~
219 255 292 0 3 22
0 52 51 50
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
3277 0 0
2
5.90019e-315 5.49149e-315
0
5 4011~
219 259 131 0 3 22
0 53 53 54
0
0 0 624 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
4212 0 0
2
5.90019e-315 5.49279e-315
0
14 Logic Display~
6 384 116 0 1 2
10 54
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.90019e-315 5.49408e-315
0
74
1 0 2 0 0 4224 0 36 0 0 35 4
826 641
693 641
693 670
688 670
2 0 3 0 0 4224 0 35 0 0 34 2
836 724
687 724
2 0 4 0 0 4096 0 36 0 0 4 4
826 659
786 659
786 699
781 699
1 3 4 0 0 4224 0 35 37 0 0 4
836 706
781 706
781 699
773 699
1 3 5 0 0 8320 0 52 23 0 0 3
1017 921
1017 931
836 931
1 3 6 0 0 8320 0 47 24 0 0 3
418 919
418 936
236 936
2 1 7 0 0 4224 0 24 7 0 0 4
185 945
133 945
133 962
124 962
1 1 8 0 0 4224 0 24 8 0 0 4
185 927
132 927
132 923
123 923
2 1 9 0 0 4224 0 23 5 0 0 4
784 940
739 940
739 958
730 958
1 1 10 0 0 4224 0 23 6 0 0 4
784 922
732 922
732 915
723 915
2 0 11 0 0 4096 0 28 0 0 12 3
719 1097
695 1097
695 1079
1 1 11 0 0 4224 0 28 2 0 0 4
719 1079
673 1079
673 1083
664 1083
2 0 12 0 0 4096 0 27 0 0 14 3
719 1166
698 1166
698 1148
1 1 12 0 0 4224 0 27 1 0 0 4
719 1148
674 1148
674 1157
665 1157
2 0 13 0 0 4096 0 32 0 0 16 3
148 1188
129 1188
129 1170
1 1 13 0 0 4224 0 32 3 0 0 4
148 1170
114 1170
114 1188
101 1188
2 0 14 0 0 8192 0 31 0 0 18 3
137 1124
122 1124
122 1106
1 1 14 0 0 4224 0 31 4 0 0 4
137 1106
111 1106
111 1109
102 1109
1 3 15 0 0 8320 0 48 25 0 0 5
1046 1113
1046 1117
999 1117
999 1111
991 1111
1 3 16 0 0 8320 0 53 29 0 0 5
430 1120
430 1144
391 1144
391 1137
383 1137
2 0 17 0 0 4096 0 25 0 0 22 3
939 1120
919 1120
919 1102
1 3 17 0 0 4224 0 25 26 0 0 4
939 1102
880 1102
880 1115
872 1115
2 0 18 0 0 4096 0 29 0 0 24 3
332 1146
313 1146
313 1128
1 3 18 0 0 4224 0 29 30 0 0 4
332 1128
289 1128
289 1139
281 1139
2 3 19 0 0 4224 0 26 27 0 0 4
820 1124
779 1124
779 1157
771 1157
1 3 20 0 0 4224 0 26 28 0 0 4
820 1106
779 1106
779 1088
771 1088
2 3 21 0 0 8320 0 30 32 0 0 4
230 1148
207 1148
207 1179
199 1179
1 3 22 0 0 4224 0 30 31 0 0 4
230 1130
196 1130
196 1115
188 1115
1 3 23 0 0 8320 0 46 33 0 0 3
1121 678
1121 681
1084 681
2 0 24 0 0 8192 0 33 0 0 31 3
1032 690
1019 690
1019 672
1 3 24 0 0 4224 0 33 34 0 0 4
1032 672
1004 672
1004 676
977 676
2 3 25 0 0 8320 0 34 35 0 0 4
925 685
911 685
911 715
888 715
1 3 26 0 0 12416 0 34 36 0 0 4
925 667
908 667
908 650
878 650
2 1 3 0 0 0 0 37 9 0 0 4
721 708
687 708
687 733
674 733
1 1 2 0 0 0 0 37 10 0 0 4
721 690
688 690
688 670
679 670
1 3 27 0 0 8320 0 50 59 0 0 3
489 733
489 745
395 745
2 3 28 0 0 4224 0 59 57 0 0 4
344 754
302 754
302 776
294 776
1 3 29 0 0 4224 0 59 60 0 0 4
344 736
301 736
301 706
293 706
1 1 30 0 0 4224 0 60 12 0 0 4
242 697
129 697
129 703
115 703
2 1 31 0 0 4224 0 57 11 0 0 4
243 785
120 785
120 776
106 776
1 0 32 0 0 4096 0 57 0 0 42 4
243 767
211 767
211 743
206 743
2 3 32 0 0 4224 0 60 58 0 0 4
242 715
206 715
206 743
198 743
2 1 31 0 0 0 0 58 11 0 0 4
147 752
115 752
115 776
106 776
1 1 30 0 0 0 0 58 12 0 0 4
147 734
124 734
124 703
115 703
2 1 33 0 0 4224 0 40 16 0 0 4
764 519
698 519
698 561
689 561
1 1 34 0 0 4224 0 40 15 0 0 4
764 501
698 501
698 481
689 481
2 0 35 0 0 4096 0 39 0 0 48 3
909 522
873 522
873 504
1 3 35 0 0 4224 0 39 40 0 0 4
909 504
824 504
824 510
816 510
1 3 36 0 0 8320 0 51 39 0 0 3
1017 501
1017 513
961 513
2 0 37 0 0 4096 0 42 0 0 53 3
726 255
706 255
706 237
2 0 38 0 0 4096 0 41 0 0 52 3
741 350
715 350
715 332
1 1 38 0 0 4224 0 41 13 0 0 4
741 332
696 332
696 345
687 345
1 1 37 0 0 4224 0 42 17 0 0 4
726 237
686 237
686 248
677 248
2 3 39 0 0 4224 0 38 41 0 0 4
911 313
801 313
801 341
793 341
1 3 40 0 0 4224 0 38 42 0 0 4
911 295
786 295
786 246
778 246
1 3 41 0 0 8320 0 44 38 0 0 3
1058 300
1058 304
963 304
2 0 42 0 0 4096 0 43 0 0 58 3
813 127
752 127
752 109
1 1 42 0 0 4224 0 43 18 0 0 4
813 109
724 109
724 125
715 125
1 3 43 0 0 8320 0 45 43 0 0 3
1020 105
1020 118
865 118
1 3 44 0 0 8320 0 49 56 0 0 3
457 522
457 529
374 529
1 3 45 0 0 4224 0 56 61 0 0 4
323 520
255 520
255 487
247 487
2 3 46 0 0 4224 0 56 55 0 0 4
323 538
258 538
258 567
250 567
2 0 47 0 0 4096 0 55 0 0 64 3
199 576
176 576
176 558
1 1 47 0 0 4224 0 55 19 0 0 4
199 558
159 558
159 575
150 575
2 0 48 0 0 4096 0 61 0 0 66 3
196 496
175 496
175 478
1 1 48 0 0 4224 0 61 14 0 0 4
196 478
161 478
161 468
152 468
1 3 49 0 0 8320 0 54 62 0 0 5
488 306
488 310
412 310
412 293
404 293
2 0 50 0 0 4096 0 62 0 0 69 3
353 302
314 302
314 284
1 3 50 0 0 4224 0 62 63 0 0 4
353 284
290 284
290 292
282 292
2 1 51 0 0 4224 0 63 20 0 0 4
231 301
187 301
187 327
178 327
1 1 52 0 0 4224 0 63 21 0 0 4
231 283
183 283
183 273
174 273
2 0 53 0 0 4096 0 64 0 0 74 3
235 140
197 140
197 122
1 3 54 0 0 8320 0 65 64 0 0 4
384 134
384 138
286 138
286 131
1 1 53 0 0 4224 0 64 22 0 0 4
235 122
179 122
179 123
170 123
159
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
219 1151 280 1175
229 1159 269 1175
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
219 1087 280 1111
229 1095 269 1111
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
316 1149 377 1173
326 1157 366 1173
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
320 1086 381 1110
330 1094 370 1110
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
379 1142 440 1166
389 1150 429 1166
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
264 1104 325 1128
274 1112 314 1128
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
181 1180 242 1204
191 1188 231 1204
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
169 1091 230 1115
179 1099 219 1115
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
104 1190 165 1214
114 1198 154 1214
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
104 1144 165 1168
114 1152 154 1168
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
91 1116 152 1140
101 1124 141 1140
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
100 1064 161 1088
110 1072 150 1088
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
237 910 298 934
247 918 287 934
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
133 939 194 963
143 947 183 963
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
130 899 191 923
140 907 180 923
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
345 754 406 778
355 762 395 778
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
341 695 402 719
351 703 391 719
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
399 717 460 741
409 725 449 741
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
271 774 332 798
281 782 321 798
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
200 763 261 787
210 771 250 787
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
203 744 264 768
213 752 253 768
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
173 720 234 744
183 728 223 744
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
106 746 167 770
116 754 156 770
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
103 727 164 751
113 735 153 751
5 (AB)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
104 709 165 733
114 717 154 733
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
275 682 336 706
285 690 325 706
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
194 690 255 714
204 698 244 714
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
196 672 257 696
206 680 246 696
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
362 502 423 526
372 510 412 526
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
279 517 340 541
289 525 329 541
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
278 498 339 522
288 506 328 522
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
250 539 311 563
260 547 300 563
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
228 461 289 485
238 469 278 485
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
153 571 214 595
163 579 203 595
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
150 530 211 554
160 538 200 554
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
145 490 206 514
155 498 195 514
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
152 446 213 470
162 454 202 470
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
413 284 474 308
423 292 463 308
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
309 296 370 320
319 304 359 320
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
307 259 368 283
317 267 357 283
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
259 291 320 315
269 299 309 315
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
182 295 243 319
192 303 232 319
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
182 259 243 283
192 267 232 283
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
292 112 353 136
302 120 342 136
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
851 1077 912 1101
861 1085 901 1101
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
990 1114 1051 1138
1000 1122 1040 1138
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
901 1122 962 1146
911 1130 951 1146
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
907 1058 968 1082
917 1066 957 1082
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
776 1120 837 1144
786 1128 826 1144
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
751 1156 812 1180
761 1164 801 1180
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
664 1164 725 1188
674 1172 714 1188
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
665 1122 726 1146
675 1130 715 1146
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
987 685 1048 709
997 693 1037 709
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
863 688 924 712
873 696 913 712
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
788 703 849 727
798 711 838 727
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
785 683 846 707
795 691 835 707
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
749 671 810 695
759 679 799 695
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
632 687 693 711
642 695 682 711
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
632 673 693 697
642 681 682 697
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
859 516 920 540
869 524 909 540
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
858 478 919 502
868 486 908 502
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
947 486 1008 510
957 494 997 510
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
772 338 833 362
782 346 822 362
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
973 278 1034 302
983 286 1023 302
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
855 306 916 330
865 314 905 330
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
857 271 918 295
867 279 907 295
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
687 305 748 329
697 313 737 329
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
672 250 733 274
682 258 722 274
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
753 122 814 146
763 130 803 146
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
750 1060 811 1084
760 1068 800 1084
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
774 1080 835 1104
784 1088 824 1104
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
663 1092 724 1116
673 1100 713 1116
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
670 1048 731 1072
680 1056 720 1072
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
828 903 889 927
838 911 878 927
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
738 940 799 964
748 948 788 964
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
732 894 793 918
742 902 782 918
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1059 651 1120 675
1069 659 1109 675
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
918 685 979 709
928 693 968 709
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
912 625 973 649
922 633 962 649
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
958 651 1019 675
968 659 1008 675
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
858 606 919 630
868 614 908 630
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
768 634 829 658
778 642 818 658
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
770 616 831 640
780 624 820 640
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
796 477 857 501
806 485 846 501
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
706 515 767 539
716 523 756 539
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
707 475 768 499
717 483 757 499
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
762 216 823 240
772 224 812 240
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
683 344 744 368
693 352 733 368
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
676 206 737 230
686 214 726 230
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
901 93 962 117
911 101 951 117
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
751 83 812 107
761 91 801 107
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
168 133 229 157
178 141 218 157
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
168 96 229 120
178 104 218 120
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1038 428 1115 452
1048 436 1104 452
7 Y=(A+B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
457 452 582 476
467 460 571 476
13 Y=(A+B)''=A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1048 214 1173 238
1058 222 1162 238
13 Y=(A.B)''=A.B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
479 237 540 261
489 245 529 261
5 Y=A.B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1033 37 1086 61
1043 45 1075 61
4 Y=A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
390 74 443 98
400 81 432 97
4 Y=A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
898 446 975 470
908 454 964 470
7 (A+B)''
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
767 442 836 466
777 450 825 466
6 (A+B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
911 247 996 271
921 255 985 271
8 (A'+B')'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
802 321 839 345
812 329 828 345
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
803 237 840 261
813 245 829 261
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
812 56 881 80
822 64 870 80
6 (A+A)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
333 473 410 497
343 481 399 497
7 (A'B')'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
231 571 268 595
241 579 257 595
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
221 431 258 455
231 439 247 455
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
372 240 449 264
382 248 438 264
7 (A.B)''
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
237 236 306 260
247 244 295 260
6 (A.B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
214 70 283 94
224 78 272 94
6 (A.A)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
605 1151 634 1175
615 1159 623 1175
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
604 1066 633 1090
614 1074 622 1090
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
44 1168 73 1192
54 1176 62 1192
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
42 1096 71 1120
52 1104 60 1120
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
661 949 690 973
671 957 679 973
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
661 900 690 924
671 908 679 924
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
70 958 99 982
80 966 88 982
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
72 902 101 926
82 910 90 926
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
620 715 649 739
630 723 638 739
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
619 658 648 682
629 666 637 682
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
46 757 75 781
56 765 64 781
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
47 689 76 713
57 697 65 713
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
625 539 654 563
635 547 643 563
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
622 470 651 494
632 478 640 494
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
88 555 117 579
98 563 106 579
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
90 456 119 480
100 464 108 480
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
624 331 653 355
634 339 642 355
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
619 234 648 258
629 242 637 258
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
120 310 149 334
130 318 138 334
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
121 259 150 283
131 267 139 283
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
651 108 680 132
661 116 669 132
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
108 111 137 135
118 119 126 135
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
87 629 300 653
97 637 289 653
24 XOR GATE USING NAND, NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
25 4 262 28
35 12 251 28
27 BASIC GATES USING NAND, NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
294 710 363 734
304 718 352 734
6 (A'+B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
295 750 364 774
305 758 353 774
6 (A+B')
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
406 741 499 765
416 749 488 765
9 (A'B+AB')
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
672 683 741 707
682 691 730 707
6 (A+B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
866 623 927 647
876 631 916 647
5 (A'B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
881 710 942 734
891 718 931 734
5 (AB')
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1011 627 1104 651
1021 635 1093 651
9 (A'B+AB')
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
301 906 370 930
311 914 359 930
6 (A.B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
371 1110 440 1134
381 1118 429 1134
6 (A+B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
884 903 953 927
894 911 942 927
6 (A+B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
977 1080 1046 1104
987 1088 1035 1104
6 (A.B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1005 608 1066 632
1015 616 1055 632
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
283 366 400 390
293 374 389 390
12  NAND TO AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
205 175 322 199
215 183 311 199
12  NAND TO NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
290 560 399 584
300 568 388 584
11  NAND TO OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
824 136 925 160
834 144 914 160
10 NOR TO NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
836 382 945 406
846 390 934 406
11  NOR TO AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
848 553 941 577
858 561 930 577
9 NOR TO OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
810 797 919 821
820 805 908 821
11  NOR TO XOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
201 828 318 852
211 836 307 852
12  NAND TO XOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
796 981 889 1005
806 989 878 1005
9  NOR GATE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
160 981 261 1005
170 989 250 1005
10  NAND GATE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
137 1231 254 1255
147 1239 243 1255
12  NAND TO NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
767 1231 884 1255
777 1239 873 1255
12  NOR TO NAND
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
