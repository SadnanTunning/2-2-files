CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1060 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
141
13 Logic Switch~
5 1059 559 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 -3 -15 5
4 Cin1
-32 16 -4 24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90019e-315 0
0
13 Logic Switch~
5 981 598 0 1 11
0 9
0
0 0 21360 90
2 0V
-4 15 10 23
2 B1
-5 28 9 36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.90019e-315 5.26354e-315
0
13 Logic Switch~
5 952 598 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 16 8 24
2 B2
-6 30 8 38
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90019e-315 5.30499e-315
0
13 Logic Switch~
5 928 598 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 15 8 23
2 B3
-6 32 8 40
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90019e-315 5.32571e-315
0
13 Logic Switch~
5 904 599 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-5 14 9 22
2 B4
-6 31 8 39
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90019e-315 5.34643e-315
0
13 Logic Switch~
5 981 400 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -27 8 -19
2 A1
-6 -43 8 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90019e-315 5.3568e-315
0
13 Logic Switch~
5 953 399 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -26 9 -18
2 A2
-3 -41 11 -33
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90019e-315 5.36716e-315
0
13 Logic Switch~
5 928 400 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 A3
-5 -42 9 -34
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90019e-315 5.37752e-315
0
13 Logic Switch~
5 902 400 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -24 6 -16
2 A4
-7 -43 7 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90019e-315 5.38788e-315
0
13 Logic Switch~
5 1929 679 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -27 8 -19
2 A8
-3 -44 11 -36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90019e-315 5.39306e-315
0
13 Logic Switch~
5 1901 679 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -26 9 -18
2 A7
-4 -43 10 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90019e-315 5.39824e-315
0
13 Logic Switch~
5 1874 679 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 A6
-5 -43 9 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90019e-315 5.40342e-315
0
13 Logic Switch~
5 1849 679 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -24 6 -16
2 A5
-5 -43 9 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90019e-315 5.4086e-315
0
13 Logic Switch~
5 2119 680 0 1 11
0 30
0
0 0 21360 270
2 0V
-7 -21 7 -13
4 Cin4
-13 -31 15 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
5.90019e-315 5.41378e-315
0
13 Logic Switch~
5 2061 678 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -27 8 -19
2 B8
-7 -44 7 -36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.90019e-315 5.41896e-315
0
13 Logic Switch~
5 2033 677 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -26 9 -18
2 B7
-3 -43 11 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.90019e-315 5.42414e-315
0
13 Logic Switch~
5 2008 678 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 B6
-5 -42 9 -34
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.90019e-315 5.42933e-315
0
13 Logic Switch~
5 1982 678 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -24 6 -16
2 B5
-7 -42 7 -34
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.90019e-315 5.43192e-315
0
13 Logic Switch~
5 189 1153 0 1 11
0 67
0
0 0 21360 270
2 0V
-8 -24 6 -16
2 B4
-7 -42 7 -34
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
317 0 0
2
5.90019e-315 5.43451e-315
0
13 Logic Switch~
5 215 1153 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 B3
-5 -42 9 -34
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3108 0 0
2
5.90019e-315 5.4371e-315
0
13 Logic Switch~
5 240 1152 0 1 11
0 69
0
0 0 21360 270
2 0V
-5 -26 9 -18
2 B2
-3 -43 11 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4299 0 0
2
5.90019e-315 5.43969e-315
0
13 Logic Switch~
5 268 1153 0 10 11
0 70 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -27 8 -19
2 B1
-7 -44 7 -36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9672 0 0
2
5.90019e-315 5.44228e-315
0
13 Logic Switch~
5 326 1155 0 1 11
0 58
0
0 0 21360 270
2 0V
-7 -21 7 -13
4 Cin3
-13 -31 15 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7876 0 0
2
5.90019e-315 5.44487e-315
0
13 Logic Switch~
5 56 1154 0 1 11
0 73
0
0 0 21360 270
2 0V
-8 -24 6 -16
2 A4
-5 -43 9 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
5.90019e-315 5.44746e-315
0
13 Logic Switch~
5 81 1154 0 10 11
0 74 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 A3
-5 -43 9 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.90019e-315 5.45005e-315
0
13 Logic Switch~
5 108 1154 0 1 11
0 75
0
0 0 21360 270
2 0V
-5 -26 9 -18
2 A2
-4 -43 10 -35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
5.90019e-315 5.45264e-315
0
13 Logic Switch~
5 136 1154 0 10 11
0 76 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -27 8 -19
2 A1
-3 -44 11 -36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
5.90019e-315 5.45523e-315
0
13 Logic Switch~
5 487 998 0 10 11
0 94 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
18 0 32 8
4 Cin2
11 -10 39 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
5.90019e-315 5.45782e-315
0
13 Logic Switch~
5 444 1005 0 1 11
0 86
0
0 0 21360 90
2 0V
-4 15 10 23
2 B1
-5 28 9 36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
5.90019e-315 5.46041e-315
0
13 Logic Switch~
5 403 1006 0 10 11
0 87 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 16 8 24
2 B2
-6 30 8 38
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
5.90019e-315 5.463e-315
0
13 Logic Switch~
5 364 1006 0 10 11
0 88 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 15 8 23
2 B3
-6 29 8 37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3409 0 0
2
5.90019e-315 5.46559e-315
0
13 Logic Switch~
5 325 1006 0 10 11
0 89 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-5 14 9 22
2 B4
-5 28 9 36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3951 0 0
2
5.90019e-315 5.46818e-315
0
13 Logic Switch~
5 407 803 0 10 11
0 98 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -27 8 -19
2 A1
-7 -46 7 -38
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
5.90019e-315 5.47077e-315
0
13 Logic Switch~
5 379 802 0 10 11
0 97 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -26 9 -18
2 A2
-7 -45 7 -37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3780 0 0
2
5.90019e-315 5.47207e-315
0
13 Logic Switch~
5 354 803 0 10 11
0 96 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 A3
-5 -45 9 -37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9265 0 0
2
5.90019e-315 5.47336e-315
0
13 Logic Switch~
5 328 803 0 10 11
0 95 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -24 6 -16
2 A4
-10 -44 4 -36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.90019e-315 5.47466e-315
0
13 Logic Switch~
5 197 570 0 1 11
0 104
0
0 0 21360 0
2 0V
-29 -3 -15 5
3 Cin
-29 16 -8 24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
5.90019e-315 5.47595e-315
0
13 Logic Switch~
5 119 609 0 1 11
0 108
0
0 0 21360 90
2 0V
-4 15 10 23
2 B1
-3 36 11 44
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.90019e-315 5.47725e-315
0
13 Logic Switch~
5 90 609 0 10 11
0 107 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 16 8 24
2 B2
-6 37 8 45
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9281 0 0
2
5.90019e-315 5.47854e-315
0
13 Logic Switch~
5 66 609 0 10 11
0 106 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 15 8 23
2 B3
-5 34 9 42
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8464 0 0
2
5.90019e-315 5.47984e-315
0
13 Logic Switch~
5 42 610 0 10 11
0 105 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-5 14 9 22
2 B4
-8 34 6 42
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7168 0 0
2
5.90019e-315 5.48113e-315
0
13 Logic Switch~
5 119 411 0 10 11
0 112 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -27 8 -19
2 A1
-7 -46 7 -38
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3171 0 0
2
5.90019e-315 5.48243e-315
0
13 Logic Switch~
5 91 410 0 10 11
0 111 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -26 9 -18
2 A2
-7 -45 7 -37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4139 0 0
2
5.90019e-315 5.48372e-315
0
13 Logic Switch~
5 66 411 0 10 11
0 110 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 A3
-5 -45 9 -37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6435 0 0
2
5.90019e-315 5.48502e-315
0
13 Logic Switch~
5 40 411 0 10 11
0 109 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -24 6 -16
2 A4
-10 -44 4 -36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5283 0 0
2
5.90019e-315 5.48631e-315
0
13 Logic Switch~
5 81 63 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-31 -1 -17 7
1 B
-50 33 -43 41
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6874 0 0
2
44606.7 0
0
13 Logic Switch~
5 78 100 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-31 -4 -17 4
1 A
-45 -39 -38 -31
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5305 0 0
2
44606.7 1
0
13 Logic Switch~
5 600 63 0 10 11
0 120 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-34 -2 -20 6
3 Cin
-58 -3 -37 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
44606.7 2
0
13 Logic Switch~
5 597 130 0 10 11
0 72 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -5 -21 3
1 A
-51 -5 -44 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
969 0 0
2
44606.7 3
0
13 Logic Switch~
5 598 97 0 10 11
0 71 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -4 -21 4
1 B
-50 -6 -43 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8402 0 0
2
44606.7 4
0
14 Logic Display~
6 1207 385 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.90019e-315 5.48761e-315
0
14 Logic Display~
6 1236 383 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
5.90019e-315 5.4889e-315
0
14 Logic Display~
6 1168 440 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.90019e-315 5.4902e-315
0
14 Logic Display~
6 1262 383 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.90019e-315 5.49149e-315
0
14 Logic Display~
6 1287 384 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
5.90019e-315 5.49279e-315
0
6 74LS83
105 1115 497 0 14 29
0 11 12 13 14 2 3 4 5 10
15 16 17 18 19
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
319 0 0
2
5.90019e-315 5.49408e-315
0
9 Inverter~
13 903 560 0 2 22
0 6 2
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U6A
781 -159 802 -151
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3976 0 0
2
5.90019e-315 5.49538e-315
0
9 Inverter~
13 927 559 0 2 22
0 7 3
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U6B
759 -157 780 -149
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
7634 0 0
2
5.90019e-315 5.49667e-315
0
9 Inverter~
13 950 559 0 2 22
0 8 4
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U6C
734 -157 755 -149
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
523 0 0
2
5.90019e-315 5.49797e-315
0
9 Inverter~
13 978 560 0 2 22
0 9 5
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U6D
707 -158 728 -150
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
6748 0 0
2
5.90019e-315 5.49926e-315
0
9 2-In XOR~
219 2216 1226 0 3 22
0 23 31 40
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U21A
1276 -239 1304 -231
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
6901 0 0
2
5.90019e-315 5.50056e-315
0
9 2-In XOR~
219 2400 1217 0 3 22
0 45 40 36
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U18D
1075 -225 1103 -217
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
842 0 0
2
5.90019e-315 5.50185e-315
0
9 2-In AND~
219 2233 1312 0 3 22
0 23 31 48
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U19C
1279 -381 1307 -373
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
3277 0 0
2
5.90019e-315 5.50315e-315
0
9 2-In AND~
219 2415 1282 0 3 22
0 40 45 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U19B
1076 -348 1104 -340
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
4212 0 0
2
5.90019e-315 5.50444e-315
0
14 Logic Display~
6 2672 664 0 1 2
10 36
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L29
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.90019e-315 5.50574e-315
0
8 2-In OR~
219 2555 1291 0 3 22
0 22 48 35
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U20A
938 -280 966 -272
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
5551 0 0
2
5.90019e-315 5.50703e-315
0
9 2-In XOR~
219 2219 1071 0 3 22
0 42 32 25
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U18C
1258 -239 1286 -231
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
6986 0 0
2
5.90019e-315 5.50833e-315
0
9 2-In XOR~
219 2415 1063 0 3 22
0 46 25 37
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U18B
1072 -297 1100 -289
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
8745 0 0
2
5.90019e-315 5.50963e-315
0
9 2-In AND~
219 2205 1155 0 3 22
0 42 32 49
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U19A
1223 -349 1251 -341
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
9592 0 0
2
5.90019e-315 5.51092e-315
0
9 2-In AND~
219 2401 1122 0 3 22
0 25 46 24
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17D
1099 -190 1127 -182
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
8748 0 0
2
5.90019e-315 5.51222e-315
0
14 Logic Display~
6 2701 665 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L28
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90019e-315 5.51286e-315
0
8 2-In OR~
219 2538 1130 0 3 22
0 24 49 45
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13D
923 -218 951 -210
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
631 0 0
2
5.90019e-315 5.51351e-315
0
9 2-In XOR~
219 2181 914 0 3 22
0 43 33 27
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U18A
1271 -4 1299 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
9466 0 0
2
5.90019e-315 5.51416e-315
0
9 2-In XOR~
219 2376 907 0 3 22
0 47 27 38
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U16D
1053 -63 1081 -55
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3266 0 0
2
5.90019e-315 5.51481e-315
0
9 2-In AND~
219 2190 1009 0 3 22
0 43 33 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17C
1259 -276 1287 -268
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
7693 0 0
2
5.90019e-315 5.51545e-315
0
9 2-In AND~
219 2377 975 0 3 22
0 27 47 41
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17B
1083 -165 1111 -157
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
3723 0 0
2
5.90019e-315 5.5161e-315
0
14 Logic Display~
6 2731 664 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L27
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
5.90019e-315 5.51675e-315
0
8 2-In OR~
219 2510 984 0 3 22
0 41 26 46
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13C
896 -111 924 -103
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
6263 0 0
2
5.90019e-315 5.5174e-315
0
8 2-In OR~
219 2485 812 0 3 22
0 28 50 47
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13B
985 -139 1013 -131
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
4900 0 0
2
5.90019e-315 5.51804e-315
0
14 Logic Display~
6 2762 665 0 1 2
10 39
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L26
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8783 0 0
2
5.90019e-315 5.51869e-315
0
9 2-In AND~
219 2336 804 0 3 22
0 30 29 28
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17A
1130 -73 1158 -65
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3221 0 0
2
5.90019e-315 5.51934e-315
0
9 2-In AND~
219 2185 848 0 3 22
0 44 34 50
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11D
1238 -51 1266 -43
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
3215 0 0
2
5.90019e-315 5.51999e-315
0
9 2-In XOR~
219 2346 741 0 3 22
0 30 29 39
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U16C
1120 140 1148 148
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
7903 0 0
2
5.90019e-315 5.52063e-315
0
9 2-In XOR~
219 2174 750 0 3 22
0 44 34 29
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U16B
1260 4 1288 12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
7121 0 0
2
5.90019e-315 5.52128e-315
0
14 Logic Display~
6 2635 665 0 1 2
10 35
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L25
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
5.90019e-315 5.52193e-315
0
14 Logic Display~
6 884 1137 0 1 2
10 53
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L24
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
5.90019e-315 5.52258e-315
0
9 2-In XOR~
219 337 1580 0 3 22
0 68 58 63
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U15B
1331 -259 1359 -251
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
7804 0 0
2
5.90019e-315 5.52322e-315
0
9 2-In XOR~
219 325 1421 0 3 22
0 69 58 65
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U15A
1354 -286 1382 -278
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
5523 0 0
2
5.90019e-315 5.52387e-315
0
9 2-In XOR~
219 321 1255 0 3 22
0 70 58 66
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12D
1351 -60 1379 -52
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
3330 0 0
2
5.90019e-315 5.52452e-315
0
9 2-In XOR~
219 322 1724 0 3 22
0 67 58 51
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U14A
1400 -646 1428 -638
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3465 0 0
2
5.90019e-315 5.52517e-315
0
6 74LS83
105 252 508 0 14 29
0 109 110 111 112 105 106 107 108 104
113 114 115 116 117
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8396 0 0
2
5.90019e-315 5.52581e-315
0
9 2-In XOR~
219 473 1224 0 3 22
0 76 66 83
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2D
1263 4 1284 12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3685 0 0
2
5.90019e-315 5.52646e-315
0
9 2-In XOR~
219 637 1215 0 3 22
0 58 83 57
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U9A
1077 108 1098 116
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7849 0 0
2
5.90019e-315 5.52711e-315
0
9 2-In AND~
219 478 1324 0 3 22
0 76 66 85
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3D
1241 -51 1262 -43
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
6343 0 0
2
5.90019e-315 5.52776e-315
0
9 2-In AND~
219 600 1281 0 3 22
0 83 58 84
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10A
1130 -73 1158 -65
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7376 0 0
2
5.90019e-315 5.52841e-315
0
14 Logic Display~
6 999 1133 0 1 2
10 57
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
5.90019e-315 5.52905e-315
0
8 2-In OR~
219 736 1290 0 3 22
0 84 85 79
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U4B
988 -139 1009 -131
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5776 0 0
2
5.90019e-315 5.5297e-315
0
8 2-In OR~
219 775 1457 0 3 22
0 64 82 78
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U4C
899 -111 920 -103
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7207 0 0
2
5.90019e-315 5.53035e-315
0
14 Logic Display~
6 971 1134 0 1 2
10 56
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L21
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
5.90019e-315 5.531e-315
0
9 2-In AND~
219 644 1448 0 3 22
0 52 79 64
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10B
1083 -165 1111 -157
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3760 0 0
2
5.90019e-315 5.53164e-315
0
9 2-In AND~
219 467 1486 0 3 22
0 75 65 82
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10C
1259 -276 1287 -268
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
754 0 0
2
5.90019e-315 5.53229e-315
0
9 2-In XOR~
219 686 1381 0 3 22
0 79 52 56
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U9B
988 -55 1009 -47
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9767 0 0
2
5.90019e-315 5.53294e-315
0
9 2-In XOR~
219 488 1390 0 3 22
0 75 65 52
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U9C
1274 -4 1295 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
7978 0 0
2
5.90019e-315 5.53359e-315
0
8 2-In OR~
219 782 1608 0 3 22
0 61 81 77
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U4D
926 -218 947 -210
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3142 0 0
2
5.90019e-315 5.53423e-315
0
14 Logic Display~
6 941 1135 0 1 2
10 55
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L22
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3284 0 0
2
5.90019e-315 5.53488e-315
0
9 2-In AND~
219 644 1599 0 3 22
0 62 78 61
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10D
1099 -190 1127 -182
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
659 0 0
2
5.90019e-315 5.53553e-315
0
9 2-In AND~
219 477 1630 0 3 22
0 74 63 81
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11A
1223 -349 1251 -341
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3800 0 0
2
5.90019e-315 5.53618e-315
0
9 2-In XOR~
219 682 1539 0 3 22
0 78 62 55
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U9D
973 -303 994 -295
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
6792 0 0
2
5.90019e-315 5.53682e-315
0
9 2-In XOR~
219 476 1548 0 3 22
0 74 63 62
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12A
1184 -237 1212 -229
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3701 0 0
2
5.90019e-315 5.53747e-315
0
8 2-In OR~
219 787 1765 0 3 22
0 59 80 53
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13A
938 -280 966 -272
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
6316 0 0
2
5.90019e-315 5.53812e-315
0
14 Logic Display~
6 912 1135 0 1 2
10 54
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L23
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8734 0 0
2
5.90019e-315 5.53877e-315
0
9 2-In AND~
219 643 1757 0 3 22
0 60 77 59
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11B
1076 -348 1104 -340
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
7988 0 0
2
5.90019e-315 5.53941e-315
0
9 2-In AND~
219 482 1787 0 3 22
0 73 51 80
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11C
1279 -381 1307 -373
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3217 0 0
2
5.90019e-315 5.54006e-315
0
9 2-In XOR~
219 646 1692 0 3 22
0 77 60 54
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12B
1075 -225 1103 -217
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3965 0 0
2
5.90019e-315 5.54071e-315
0
9 2-In XOR~
219 475 1701 0 3 22
0 73 51 60
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12C
1276 -239 1304 -231
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
8239 0 0
2
5.90019e-315 5.54136e-315
0
9 2-In XOR~
219 433 956 0 3 22
0 94 86 93
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U7D
-429 -123 -408 -115
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
828 0 0
2
5.90019e-315 5.542e-315
0
9 2-In XOR~
219 392 952 0 3 22
0 94 87 92
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U7C
-386 -129 -365 -121
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6187 0 0
2
5.90019e-315 5.54265e-315
0
9 2-In XOR~
219 353 956 0 3 22
0 94 88 91
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U7B
-347 -145 -326 -137
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7107 0 0
2
5.90019e-315 5.5433e-315
0
9 2-In XOR~
219 314 957 0 3 22
0 94 89 90
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U7A
-306 -161 -285 -153
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6433 0 0
2
5.90019e-315 5.54395e-315
0
14 Logic Display~
6 633 788 0 1 2
10 99
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8559 0 0
2
5.90019e-315 5.54459e-315
0
14 Logic Display~
6 662 786 0 1 2
10 100
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3674 0 0
2
5.90019e-315 5.54524e-315
0
14 Logic Display~
6 600 789 0 1 2
10 103
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5697 0 0
2
5.90019e-315 5.54589e-315
0
14 Logic Display~
6 688 786 0 1 2
10 101
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3805 0 0
2
5.90019e-315 5.54654e-315
0
14 Logic Display~
6 713 787 0 1 2
10 102
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5219 0 0
2
5.90019e-315 5.54719e-315
0
6 74LS83
105 541 900 0 14 29
0 95 96 97 98 90 91 92 93 94
99 100 101 102 103
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3795 0 0
2
5.90019e-315 5.54783e-315
0
14 Logic Display~
6 345 396 0 1 2
10 113
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3637 0 0
2
5.90019e-315 5.54848e-315
0
14 Logic Display~
6 374 394 0 1 2
10 114
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
5.90019e-315 5.54913e-315
0
14 Logic Display~
6 316 395 0 1 2
10 117
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6966 0 0
2
5.90019e-315 5.54978e-315
0
14 Logic Display~
6 400 394 0 1 2
10 115
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9796 0 0
2
5.90019e-315 5.55042e-315
0
14 Logic Display~
6 425 395 0 1 2
10 116
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5952 0 0
2
5.90019e-315 5.55107e-315
0
9 2-In XOR~
219 196 80 0 3 22
0 21 20 118
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3649 0 0
2
44606.7 5
0
9 2-In AND~
219 213 181 0 3 22
0 21 20 119
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3716 0 0
2
44606.7 6
0
14 Logic Display~
6 280 76 0 1 2
10 118
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L6
-10 -11 4 -3
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
44606.7 7
0
14 Logic Display~
6 284 177 0 1 2
10 119
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L7
-11 -15 3 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4681 0 0
2
44606.7 8
0
9 2-In XOR~
219 749 106 0 3 22
0 71 72 121
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9730 0 0
2
44606.7 9
0
9 2-In XOR~
219 941 97 0 3 22
0 120 121 122
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9874 0 0
2
44606.7 10
0
9 2-In AND~
219 773 225 0 3 22
0 72 71 125
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3B
-13 -27 8 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
364 0 0
2
44606.7 11
0
9 2-In AND~
219 932 181 0 3 22
0 121 120 124
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3656 0 0
2
44606.7 12
0
14 Logic Display~
6 1202 92 0 1 2
10 122
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3131 0 0
2
44606.7 13
0
14 Logic Display~
6 1202 186 0 1 2
10 123
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L9
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6772 0 0
2
44606.7 14
0
8 2-In OR~
219 1067 190 0 3 22
0 124 125 123
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9557 0 0
2
44606.7 15
0
170
2 5 2 0 0 8320 0 57 56 0 0 3
906 542
906 497
1083 497
2 6 3 0 0 8320 0 58 56 0 0 3
930 541
930 506
1083 506
2 7 4 0 0 8320 0 59 56 0 0 3
953 541
953 515
1083 515
2 8 5 0 0 8320 0 60 56 0 0 3
981 542
981 524
1083 524
1 1 6 0 0 4224 0 57 5 0 0 3
906 578
906 586
905 586
1 1 7 0 0 4224 0 58 4 0 0 3
930 577
930 585
929 585
1 1 8 0 0 4224 0 59 3 0 0 2
953 577
953 585
1 1 9 0 0 4224 0 60 2 0 0 3
981 578
981 585
982 585
1 9 10 0 0 8320 0 1 56 0 0 4
1071 559
1080 559
1080 542
1083 542
1 1 11 0 0 8320 0 9 56 0 0 3
902 412
902 461
1083 461
1 2 12 0 0 8320 0 8 56 0 0 3
928 412
928 470
1083 470
1 3 13 0 0 8320 0 7 56 0 0 3
953 411
953 479
1083 479
1 4 14 0 0 8320 0 6 56 0 0 3
981 412
981 488
1083 488
10 1 15 0 0 8320 0 56 51 0 0 3
1147 488
1207 488
1207 403
11 1 16 0 0 8320 0 56 52 0 0 3
1147 497
1236 497
1236 401
12 1 17 0 0 4224 0 56 54 0 0 3
1147 506
1262 506
1262 401
13 1 18 0 0 4224 0 56 55 0 0 3
1147 515
1287 515
1287 402
14 1 19 0 0 8320 0 56 53 0 0 3
1147 542
1168 542
1168 458
2 0 20 0 0 8320 0 132 0 0 21 4
189 190
104 190
104 100
99 100
1 0 21 0 0 8320 0 132 0 0 162 3
189 172
142 172
142 63
2 1 20 0 0 0 0 131 47 0 0 4
180 89
99 89
99 100
90 100
3 1 22 0 0 4224 0 64 66 0 0 2
2436 1282
2542 1282
1 0 23 0 0 8192 0 63 0 0 48 3
2209 1303
2128 1303
2128 1218
3 1 24 0 0 4224 0 70 72 0 0 4
2422 1122
2517 1122
2517 1121
2525 1121
1 0 25 0 0 4096 0 70 0 0 63 3
2377 1113
2320 1113
2320 1071
2 3 26 0 0 12416 0 78 75 0 0 4
2497 993
2393 993
2393 1009
2211 1009
1 0 27 0 0 4096 0 76 0 0 28 3
2353 966
2283 966
2283 914
3 2 27 0 0 4224 0 73 74 0 0 4
2214 914
2352 914
2352 916
2360 916
3 1 28 0 0 4224 0 81 79 0 0 4
2357 804
2464 804
2464 803
2472 803
2 0 29 0 0 4096 0 81 0 0 66 3
2312 813
2238 813
2238 750
1 0 30 0 0 8192 0 81 0 0 45 3
2312 795
2255 795
2255 732
2 0 31 0 0 4096 0 63 0 0 33 3
2209 1321
2100 1321
2100 1235
1 2 31 0 0 4224 0 18 61 0 0 3
1982 690
1982 1235
2200 1235
2 0 32 0 0 4096 0 69 0 0 35 3
2181 1164
2091 1164
2091 1082
1 2 32 0 0 4224 0 17 67 0 0 5
2008 690
2008 1082
2091 1082
2091 1080
2203 1080
2 0 33 0 0 8192 0 75 0 0 37 3
2166 1018
2087 1018
2087 924
1 2 33 0 0 4224 0 16 73 0 0 5
2033 689
2033 924
2087 924
2087 923
2165 923
2 0 34 0 0 8320 0 82 0 0 39 3
2161 857
2084 857
2084 758
1 2 34 0 0 0 0 15 84 0 0 5
2061 690
2061 758
2084 758
2084 759
2158 759
3 1 35 0 0 8320 0 66 85 0 0 3
2588 1291
2635 1291
2635 683
3 1 36 0 0 8320 0 62 65 0 0 3
2433 1217
2672 1217
2672 682
3 1 37 0 0 8320 0 68 71 0 0 3
2448 1063
2701 1063
2701 683
3 1 38 0 0 4224 0 74 77 0 0 4
2409 907
2732 907
2732 682
2731 682
3 1 39 0 0 4224 0 83 80 0 0 3
2379 741
2762 741
2762 683
1 1 30 0 0 12416 0 14 83 0 0 6
2119 692
2120 692
2120 708
2255 708
2255 732
2330 732
1 0 40 0 0 4096 0 64 0 0 60 3
2391 1273
2321 1273
2321 1226
3 1 41 0 0 4224 0 76 78 0 0 2
2398 975
2497 975
1 1 23 0 0 16512 0 61 13 0 0 5
2200 1217
2190 1217
2190 1218
1849 1218
1849 691
1 0 42 0 0 8192 0 69 0 0 50 3
2181 1146
2118 1146
2118 1064
1 1 42 0 0 16512 0 67 12 0 0 5
2203 1062
2118 1062
2118 1064
1874 1064
1874 691
1 0 43 0 0 8192 0 75 0 0 52 3
2166 1000
2108 1000
2108 906
1 1 43 0 0 16512 0 73 11 0 0 5
2165 905
2108 905
2108 906
1901 906
1901 691
1 0 44 0 0 8192 0 82 0 0 54 3
2161 839
2103 839
2103 740
1 1 44 0 0 8320 0 10 84 0 0 5
1929 691
1929 740
2103 740
2103 741
2158 741
0 1 45 0 0 4096 0 0 62 58 0 2
2305 1208
2384 1208
1 0 46 0 0 4096 0 68 0 0 61 4
2399 1054
2317 1054
2317 1055
2302 1055
1 0 47 0 0 4096 0 74 0 0 64 4
2360 898
2280 898
2280 897
2265 897
2 3 45 0 0 12416 0 64 72 0 0 6
2391 1291
2305 1291
2305 1177
2580 1177
2580 1130
2571 1130
3 2 48 0 0 4224 0 63 66 0 0 4
2254 1312
2439 1312
2439 1300
2542 1300
3 2 40 0 0 4224 0 61 62 0 0 2
2249 1226
2384 1226
2 3 46 0 0 12416 0 70 78 0 0 6
2377 1131
2302 1131
2302 1030
2552 1030
2552 984
2543 984
3 2 49 0 0 4224 0 69 72 0 0 4
2226 1155
2421 1155
2421 1139
2525 1139
3 2 25 0 0 4224 0 67 68 0 0 3
2252 1071
2399 1071
2399 1072
2 3 47 0 0 12416 0 76 79 0 0 6
2353 984
2265 984
2265 861
2523 861
2523 812
2518 812
3 2 50 0 0 4224 0 82 79 0 0 4
2206 848
2355 848
2355 821
2472 821
3 2 29 0 0 4224 0 84 83 0 0 2
2207 750
2330 750
2 0 51 0 0 4224 0 113 0 0 68 3
458 1796
369 1796
369 1724
3 2 51 0 0 0 0 90 115 0 0 4
355 1724
385 1724
385 1710
459 1710
1 0 52 0 0 8192 0 100 0 0 70 3
620 1439
573 1439
573 1390
3 2 52 0 0 4224 0 103 102 0 0 2
521 1390
670 1390
3 1 53 0 0 8320 0 110 86 0 0 3
820 1765
884 1765
884 1155
3 1 54 0 0 8320 0 114 111 0 0 3
679 1692
912 1692
912 1153
3 1 55 0 0 8320 0 108 105 0 0 3
715 1539
941 1539
941 1153
3 1 56 0 0 4224 0 102 99 0 0 4
719 1381
970 1381
970 1152
971 1152
3 1 57 0 0 4224 0 93 96 0 0 3
670 1215
999 1215
999 1151
2 0 58 0 0 4096 0 87 0 0 79 2
321 1589
284 1589
2 0 58 0 0 0 0 88 0 0 79 2
309 1430
284 1430
2 0 58 0 0 0 0 89 0 0 79 2
305 1264
284 1264
1 2 58 0 0 12416 0 23 90 0 0 5
326 1167
326 1170
284 1170
284 1733
306 1733
1 1 58 0 0 0 0 23 93 0 0 6
326 1167
327 1167
327 1170
564 1170
564 1206
621 1206
1 3 59 0 0 12416 0 110 112 0 0 4
774 1756
771 1756
771 1757
664 1757
1 0 60 0 0 4096 0 112 0 0 114 3
619 1748
563 1748
563 1701
1 3 61 0 0 4224 0 104 106 0 0 2
769 1599
665 1599
1 0 62 0 0 4096 0 106 0 0 117 3
620 1590
567 1590
567 1548
0 2 63 0 0 8320 0 0 107 90 0 3
375 1580
375 1639
453 1639
3 1 64 0 0 4224 0 100 98 0 0 2
665 1448
762 1448
2 0 65 0 0 4224 0 101 0 0 91 4
443 1495
362 1495
362 1422
361 1422
0 2 66 0 0 4224 0 0 94 92 0 3
377 1233
377 1333
454 1333
2 0 58 0 0 0 0 95 0 0 80 3
576 1290
511 1290
511 1170
3 2 63 0 0 0 0 87 109 0 0 4
370 1580
387 1580
387 1557
460 1557
3 2 65 0 0 0 0 88 103 0 0 6
358 1421
361 1421
361 1422
396 1422
396 1399
472 1399
3 2 66 0 0 0 0 89 92 0 0 4
354 1255
362 1255
362 1233
457 1233
1 1 67 0 0 4224 0 19 90 0 0 3
189 1165
189 1715
306 1715
1 1 68 0 0 4224 0 20 87 0 0 3
215 1165
215 1571
321 1571
1 1 69 0 0 4224 0 21 88 0 0 3
240 1164
240 1412
309 1412
1 1 70 0 0 4224 0 22 89 0 0 3
268 1165
268 1246
305 1246
2 0 71 0 0 8320 0 137 0 0 99 3
749 234
655 234
655 97
1 0 72 0 0 8320 0 137 0 0 100 3
749 216
676 216
676 130
1 1 71 0 0 0 0 50 135 0 0 2
610 97
733 97
1 2 72 0 0 0 0 49 135 0 0 4
609 130
692 130
692 115
733 115
1 0 73 0 0 8192 0 113 0 0 102 4
458 1778
396 1778
396 1693
397 1693
1 1 73 0 0 16512 0 115 24 0 0 5
459 1692
397 1692
397 1693
56 1693
56 1166
1 0 74 0 0 8192 0 107 0 0 104 3
453 1621
396 1621
396 1539
1 1 74 0 0 4224 0 109 25 0 0 3
460 1539
81 1539
81 1166
1 0 75 0 0 8192 0 101 0 0 106 3
443 1477
383 1477
383 1381
1 1 75 0 0 4224 0 103 26 0 0 3
472 1381
108 1381
108 1166
1 0 76 0 0 8192 0 94 0 0 108 3
454 1315
397 1315
397 1215
1 1 76 0 0 8320 0 27 92 0 0 3
136 1166
136 1215
457 1215
0 1 77 0 0 4096 0 0 114 112 0 2
551 1683
630 1683
1 0 78 0 0 4096 0 108 0 0 115 2
666 1530
555 1530
1 0 79 0 0 4096 0 102 0 0 118 2
670 1372
561 1372
2 3 77 0 0 12416 0 112 104 0 0 6
619 1766
551 1766
551 1652
822 1652
822 1608
815 1608
3 2 80 0 0 4224 0 113 110 0 0 4
503 1787
665 1787
665 1774
774 1774
3 2 60 0 0 4224 0 115 114 0 0 2
508 1701
630 1701
2 3 78 0 0 12416 0 106 98 0 0 6
620 1608
555 1608
555 1505
816 1505
816 1457
808 1457
3 2 81 0 0 4224 0 107 104 0 0 4
498 1630
660 1630
660 1617
769 1617
3 2 62 0 0 4224 0 109 108 0 0 2
509 1548
666 1548
2 3 79 0 0 12416 0 100 97 0 0 6
620 1457
561 1457
561 1336
787 1336
787 1290
769 1290
3 2 82 0 0 4224 0 101 98 0 0 4
488 1486
665 1486
665 1466
762 1466
1 0 83 0 0 8192 0 95 0 0 123 3
576 1272
530 1272
530 1224
3 1 84 0 0 4224 0 95 97 0 0 2
621 1281
723 1281
3 2 85 0 0 4224 0 94 97 0 0 4
499 1324
620 1324
620 1299
723 1299
3 2 83 0 0 4224 0 92 93 0 0 2
506 1224
621 1224
2 1 86 0 0 4224 0 116 29 0 0 2
445 975
445 992
2 1 87 0 0 4224 0 117 30 0 0 2
404 971
404 993
2 1 88 0 0 4224 0 118 31 0 0 2
365 975
365 993
2 1 89 0 0 4224 0 119 32 0 0 2
326 976
326 993
3 5 90 0 0 8320 0 119 125 0 0 3
317 927
317 900
509 900
3 6 91 0 0 8320 0 118 125 0 0 3
356 926
356 909
509 909
3 7 92 0 0 8320 0 117 125 0 0 3
395 922
395 918
509 918
3 8 93 0 0 4224 0 116 125 0 0 4
436 926
501 926
501 927
509 927
1 0 94 0 0 4096 0 116 0 0 135 2
427 975
427 985
1 0 94 0 0 4096 0 117 0 0 135 2
386 971
386 985
1 0 94 0 0 0 0 118 0 0 135 3
347 975
347 985
345 985
1 1 94 0 0 4224 0 28 119 0 0 3
488 985
308 985
308 976
9 1 94 0 0 0 0 125 28 0 0 3
509 945
488 945
488 985
1 1 95 0 0 8320 0 36 125 0 0 3
328 815
328 864
509 864
1 2 96 0 0 8320 0 35 125 0 0 3
354 815
354 873
509 873
1 3 97 0 0 8320 0 34 125 0 0 3
379 814
379 882
509 882
1 4 98 0 0 8320 0 33 125 0 0 3
407 815
407 891
509 891
10 1 99 0 0 8320 0 125 120 0 0 3
573 891
633 891
633 806
11 1 100 0 0 8320 0 125 121 0 0 3
573 900
662 900
662 804
12 1 101 0 0 4224 0 125 123 0 0 3
573 909
688 909
688 804
13 1 102 0 0 4224 0 125 124 0 0 3
573 918
713 918
713 805
14 1 103 0 0 8320 0 125 122 0 0 3
573 945
600 945
600 807
1 9 104 0 0 8320 0 37 91 0 0 4
209 570
218 570
218 553
220 553
1 5 105 0 0 8320 0 41 91 0 0 3
43 597
43 508
220 508
1 6 106 0 0 8320 0 40 91 0 0 3
67 596
67 517
220 517
1 7 107 0 0 8320 0 39 91 0 0 3
91 596
91 526
220 526
1 8 108 0 0 8320 0 38 91 0 0 3
120 596
120 535
220 535
1 1 109 0 0 8320 0 45 91 0 0 3
40 423
40 472
220 472
1 2 110 0 0 8320 0 44 91 0 0 3
66 423
66 481
220 481
1 3 111 0 0 8320 0 43 91 0 0 3
91 422
91 490
220 490
1 4 112 0 0 8320 0 42 91 0 0 3
119 423
119 499
220 499
10 1 113 0 0 8320 0 91 126 0 0 3
284 499
345 499
345 414
11 1 114 0 0 8320 0 91 127 0 0 3
284 508
374 508
374 412
12 1 115 0 0 4224 0 91 129 0 0 3
284 517
400 517
400 412
13 1 116 0 0 4224 0 91 130 0 0 3
284 526
425 526
425 413
14 1 117 0 0 8320 0 91 128 0 0 3
284 553
316 553
316 413
1 3 118 0 0 4224 0 133 131 0 0 2
264 80
229 80
1 3 119 0 0 4224 0 134 132 0 0 2
268 181
234 181
1 1 21 0 0 0 0 46 131 0 0 4
93 63
172 63
172 71
180 71
2 0 120 0 0 8192 0 138 0 0 169 3
908 190
834 190
834 88
1 0 121 0 0 8192 0 138 0 0 170 3
908 172
854 172
854 106
1 3 122 0 0 4224 0 139 136 0 0 4
1186 96
989 96
989 97
974 97
1 3 123 0 0 4224 0 140 141 0 0 2
1186 190
1100 190
3 1 124 0 0 4224 0 138 141 0 0 2
953 181
1054 181
3 2 125 0 0 4224 0 137 141 0 0 4
794 225
942 225
942 199
1054 199
1 1 120 0 0 4224 0 48 136 0 0 4
612 63
779 63
779 88
925 88
3 2 121 0 0 4224 0 135 136 0 0 2
782 106
925 106
90
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1120 386 1208 409
1132 396 1195 411
9 CARRY BIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1083 167 1145 190
1096 177 1131 192
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1004 191 1064 214
1016 201 1051 216
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
998 159 1060 182
1011 169 1046 184
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
937 151 997 174
949 161 984 176
5 PIN-6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
857 182 919 205
870 192 905 207
5 PIN-5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
858 141 920 164
871 151 906 166
5 PIN-4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
963 67 1023 90
975 77 1010 92
5 PIN-6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
875 100 935 123
887 110 922 125
5 PIN-5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
876 59 938 82
889 69 924 84
5 PIN-4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
766 100 828 123
779 110 814 125
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
778 220 840 243
791 230 826 245
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
703 226 763 249
715 236 750 251
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
698 189 760 212
711 199 746 214
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
685 108 745 131
697 118 732 133
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
672 70 734 93
685 80 720 95
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
212 53 274 76
225 63 260 78
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
143 184 203 207
155 194 190 209
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
141 144 203 167
154 154 189 169
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
218 174 280 197
231 184 266 199
5 PIN-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
134 81 194 104
146 91 181 106
5 PIN-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
122 34 184 57
135 44 170 59
5 PIN-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
565 968 705 991
578 978 691 993
16 ADDER+SUBTRACTOR
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2327 1183 2386 1206
2335 1190 2377 1205
6 Pin-12
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2328 1225 2387 1248
2336 1233 2378 1248
6 Pin-13
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2435 1192 2494 1215
2443 1199 2485 1214
6 Pin-11
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2143 1232 2202 1255
2151 1239 2193 1254
6 Pin-10
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2140 1193 2192 1216
2148 1200 2183 1215
5 Pin-9
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2244 1225 2298 1248
2253 1232 2288 1247
5 Pin-8
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2424 1252 2483 1275
2432 1259 2474 1274
6 Pin-11
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2328 1250 2387 1273
2336 1257 2378 1272
6 Pin-12
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2335 1286 2394 1309
2343 1294 2385 1309
6 Pin-13
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2152 1276 2211 1299
2160 1283 2202 1298
6 Pin-10
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2253 1312 2305 1335
2261 1320 2296 1335
5 Pin-8
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2142 1320 2194 1343
2150 1327 2185 1342
5 Pin-9
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2289 978 2348 1001
2297 986 2339 1001
6 Pin-13
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2291 941 2350 964
2299 948 2341 963
6 Pin-12
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2387 951 2446 974
2395 958 2437 973
6 Pin-11
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2110 974 2171 997
2119 982 2161 997
6 Pin-10
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2111 1015 2163 1038
2119 1022 2154 1037
5 Pin-9
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2204 985 2256 1008
2212 992 2247 1007
5 Pin-8
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2584 1266 2643 1289
2592 1273 2634 1288
6 Pin-11
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2479 1293 2538 1316
2487 1301 2529 1316
6 Pin-13
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2484 1259 2543 1282
2492 1266 2534 1281
6 Pin-12
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2467 1138 2528 1161
2476 1145 2518 1160
6 Pin-10
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2480 1094 2534 1117
2489 1102 2524 1117
5 Pin-9
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2578 1141 2630 1164
2586 1148 2621 1163
5 Pin-8
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2550 989 2604 1012
2559 997 2594 1012
5 Pin-6
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2448 989 2500 1012
2456 996 2491 1011
5 Pin-5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2451 951 2503 974
2459 958 2494 973
5 Pin-4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2347 778 2399 801
2355 785 2390 800
5 Pin-6
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2262 808 2314 831
2270 815 2305 830
5 Pin-5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2259 771 2311 794
2267 778 2302 793
5 Pin-4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2109 854 2163 877
2118 861 2153 876
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2524 824 2576 847
2532 831 2567 846
5 Pin-3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2404 818 2458 841
2413 825 2448 840
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2412 777 2466 800
2421 784 2456 799
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2113 815 2167 838
2122 822 2157 837
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2127 1120 2181 1143
2136 1127 2171 1142
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2128 1163 2182 1186
2137 1170 2172 1185
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2218 1130 2270 1153
2226 1137 2261 1152
5 Pin-3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2332 1092 2384 1115
2340 1099 2375 1114
5 Pin-4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2336 1126 2388 1149
2344 1133 2379 1148
5 Pin-5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2413 1094 2465 1117
2421 1101 2456 1116
5 Pin-6
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2108 713 2162 736
2117 720 2152 735
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2109 757 2163 780
2118 764 2153 779
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2198 722 2252 743
2207 730 2242 745
5 Pin-3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2271 706 2323 729
2279 713 2314 728
5 Pin-4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2270 747 2324 768
2279 755 2314 770
5 Pin-5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2378 714 2432 735
2387 722 2422 737
5 Pin-6
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2205 915 2259 938
2214 922 2249 937
5 Pin-8
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2113 881 2167 904
2122 889 2157 904
5 Pin-9
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2111 920 2172 943
2120 927 2162 942
6 Pin-10
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2408 879 2467 902
2416 886 2458 901
6 Pin-11
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2290 872 2349 895
2298 879 2340 894
6 Pin-12
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
2293 910 2352 933
2301 918 2343 933
6 Pin-13
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2137 1039 2191 1060
2146 1047 2181 1062
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2140 1077 2194 1098
2149 1085 2184 1100
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2242 1047 2296 1068
2251 1055 2286 1070
5 Pin-3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2334 1032 2386 1055
2342 1039 2377 1054
5 Pin-4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2334 1067 2386 1090
2342 1074 2377 1089
5 Pin-5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
2439 1037 2493 1058
2448 1045 2483 1060
5 Pin-6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
186 219 283 242
199 229 269 244
10 HALF ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
307 57 355 80
320 67 341 82
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
305 166 365 189
317 176 352 191
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
900 251 995 274
912 261 982 276
10 FULL ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1234 72 1280 95
1246 82 1267 97
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1231 170 1293 193
1244 180 1279 195
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
235 597 400 620
247 607 387 622
20 4-BIT PARALLEL ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1138 584 1235 607
1151 594 1221 609
10 SUBTRACTOR
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
