CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
170 890 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
76 E:\2.2 - Study materials\CSE 210 (Digital Logic & System Design LAB)\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 811 168 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90021e-315 0
0
13 Logic Switch~
5 414 599 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90021e-315 5.26354e-315
0
13 Logic Switch~
5 417 801 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90021e-315 5.30499e-315
0
13 Logic Switch~
5 533 581 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90021e-315 5.32571e-315
0
13 Logic Switch~
5 535 877 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90021e-315 5.34643e-315
0
13 Logic Switch~
5 244 1018 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90021e-315 5.3568e-315
0
13 Logic Switch~
5 232 1125 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90021e-315 5.36716e-315
0
13 Logic Switch~
5 638 981 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90021e-315 5.37752e-315
0
13 Logic Switch~
5 637 1334 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90021e-315 5.38788e-315
0
13 Logic Switch~
5 324 344 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
44619.8 0
0
13 Logic Switch~
5 324 130 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
44619.8 1
0
13 Logic Switch~
5 231 238 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
44619.8 2
0
5 4011~
219 1021 177 0 3 22
0 3 8 7
0
0 0 608 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 3 0
1 U
3536 0 0
2
5.90021e-315 5.39306e-315
0
5 4011~
219 1023 294 0 3 22
0 8 2 6
0
0 0 608 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 3 0
1 U
4597 0 0
2
5.90021e-315 5.39824e-315
0
5 4011~
219 1208 186 0 3 22
0 7 5 4
0
0 0 608 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 3 0
1 U
3835 0 0
2
5.90021e-315 5.40342e-315
0
5 4011~
219 1217 285 0 3 22
0 4 6 5
0
0 0 608 0
4 4011
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 3 0
1 U
3670 0 0
2
5.90021e-315 5.4086e-315
0
7 Pulser~
4 922 240 0 10 12
0 8 33 8 34 0 0 5 5 4
7
0
0 0 4640 0
0
3 CLK
-10 -35 11 -27
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5616 0 0
2
5.90021e-315 5.41378e-315
0
14 Logic Display~
6 1370 154 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90021e-315 5.41896e-315
0
14 Logic Display~
6 1377 254 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90021e-315 5.42414e-315
0
9 Inverter~
13 828 223 0 2 22
0 3 2
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 NOT
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3108 0 0
2
5.90021e-315 5.42933e-315
0
6 74112~
219 564 726 0 7 32
0 15 12 13 11 14 9 10
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
4299 0 0
2
5.90021e-315 5.43192e-315
0
7 Pulser~
4 413 713 0 10 12
0 13 35 13 36 0 0 5 5 4
7
0
0 0 4640 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9672 0 0
2
5.90021e-315 5.43451e-315
0
14 Logic Display~
6 643 658 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.90021e-315 5.4371e-315
0
14 Logic Display~
6 671 690 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.90021e-315 5.43969e-315
0
9 2-In AND~
219 381 1069 0 3 22
0 26 17 23
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9172 0 0
2
5.90021e-315 5.44228e-315
0
9 2-In AND~
219 388 1189 0 3 22
0 24 16 22
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
7100 0 0
2
5.90021e-315 5.44487e-315
0
9 Inverter~
13 247 1156 0 2 22
0 25 24
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 NOT
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
3820 0 0
2
5.90021e-315 5.44746e-315
0
8 2-In OR~
219 499 1126 0 3 22
0 23 22 19
0
0 0 608 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7678 0 0
2
5.90021e-315 5.45005e-315
0
5 7474~
219 692 1162 0 6 22
0 21 19 18 20 17 16
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 1 0
1 U
961 0 0
2
5.90021e-315 5.45264e-315
0
7 Pulser~
4 614 1179 0 10 12
0 18 37 18 38 0 0 5 5 4
7
0
0 0 4640 0
0
3 CLK
-11 -35 10 -27
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3178 0 0
2
5.90021e-315 5.45523e-315
0
14 Logic Display~
6 845 1095 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90021e-315 5.45782e-315
0
14 Logic Display~
6 881 1117 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.90021e-315 5.46041e-315
0
14 Logic Display~
6 529 234 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
44619.8 3
0
14 Logic Display~
6 499 220 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
44619.8 4
0
7 Pulser~
4 248 288 0 10 12
0 29 39 29 40 0 0 5 5 4
7
0
0 0 4640 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9265 0 0
2
44619.8 5
0
5 7474~
219 397 274 0 6 22
0 28 30 29 27 31 32
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U1A
20 -61 41 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 1 0
1 U
9442 0 0
2
44619.8 6
0
41
2 2 2 0 0 8320 0 20 14 0 0 3
831 241
831 303
999 303
1 0 3 0 0 4096 0 20 0 0 9 2
831 205
831 168
1 0 4 0 0 12416 0 16 0 0 6 5
1193 276
1135 276
1135 249
1290 249
1290 186
2 0 5 0 0 12416 0 15 0 0 5 5
1184 195
1135 195
1135 234
1304 234
1304 285
1 3 5 0 0 0 0 19 16 0 0 3
1377 272
1377 285
1244 285
3 1 4 0 0 0 0 15 18 0 0 3
1235 186
1370 186
1370 172
3 2 6 0 0 4224 0 14 16 0 0 2
1050 294
1193 294
3 1 7 0 0 4224 0 13 15 0 0 2
1048 177
1184 177
1 1 3 0 0 4224 0 1 13 0 0 2
823 168
997 168
1 0 8 0 0 8192 0 14 0 0 12 3
999 285
960 285
960 230
0 2 8 0 0 0 0 0 13 12 0 3
960 217
960 186
997 186
1 3 8 0 0 12416 0 17 17 0 0 6
898 231
888 231
888 217
960 217
960 231
946 231
1 6 9 0 0 4224 0 24 21 0 0 4
671 708
593 708
593 708
594 708
1 7 10 0 0 8320 0 23 21 0 0 3
643 676
643 690
588 690
1 4 11 0 0 4224 0 3 21 0 0 4
429 801
526 801
526 708
540 708
1 2 12 0 0 4224 0 2 21 0 0 4
426 599
526 599
526 690
540 690
3 0 13 0 0 4224 0 21 0 0 18 2
534 699
450 699
1 3 13 0 0 0 0 22 22 0 0 6
389 704
378 704
378 679
450 679
450 704
437 704
1 5 14 0 0 8320 0 5 21 0 0 3
547 877
564 877
564 738
1 1 15 0 0 8320 0 4 21 0 0 3
545 581
564 581
564 663
2 0 16 0 0 12416 0 26 0 0 24 5
364 1198
310 1198
310 1259
759 1259
759 1126
2 0 17 0 0 12416 0 25 0 0 23 5
357 1078
310 1078
310 1025
772 1025
772 1144
1 5 17 0 0 0 0 32 29 0 0 3
881 1135
881 1144
722 1144
1 6 16 0 0 0 0 31 29 0 0 5
845 1113
845 1126
715 1126
715 1126
716 1126
0 3 18 0 0 8192 0 0 29 26 0 3
643 1156
643 1144
668 1144
1 3 18 0 0 12416 0 30 30 0 0 6
590 1170
580 1170
580 1156
652 1156
652 1170
638 1170
3 2 19 0 0 4224 0 28 29 0 0 2
532 1126
668 1126
1 4 20 0 0 8320 0 9 29 0 0 3
649 1334
692 1334
692 1174
1 1 21 0 0 8320 0 8 29 0 0 3
650 981
692 981
692 1099
3 2 22 0 0 4224 0 26 28 0 0 4
409 1189
478 1189
478 1135
486 1135
3 1 23 0 0 4224 0 25 28 0 0 4
402 1069
478 1069
478 1117
486 1117
2 1 24 0 0 8320 0 27 26 0 0 3
250 1174
250 1180
364 1180
1 1 25 0 0 8320 0 7 27 0 0 5
244 1125
249 1125
249 1136
250 1136
250 1138
1 1 26 0 0 8320 0 6 25 0 0 3
256 1018
256 1060
357 1060
1 4 27 0 0 4224 0 10 36 0 0 4
336 344
396 344
396 286
397 286
1 1 28 0 0 8320 0 11 36 0 0 3
336 130
397 130
397 211
0 3 29 0 0 4224 0 0 36 38 0 4
286 263
365 263
365 256
373 256
1 3 29 0 0 0 0 35 35 0 0 6
224 279
214 279
214 258
286 258
286 279
272 279
1 2 30 0 0 4224 0 12 36 0 0 2
243 238
373 238
1 5 31 0 0 8320 0 33 36 0 0 3
529 252
529 256
427 256
1 6 32 0 0 4224 0 34 36 0 0 4
499 238
420 238
420 238
421 238
41
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
390 1044 417 1066
399 1051 407 1067
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
344 1075 371 1097
353 1083 361 1099
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
344 1030 371 1052
353 1037 361 1053
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
229 1152 256 1174
238 1159 246 1175
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
228 1119 255 1141
237 1126 245 1142
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1036 152 1063 174
1045 159 1053 175
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
970 181 997 203
979 188 987 204
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
970 142 997 164
979 149 987 165
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
809 223 838 245
819 231 827 247
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
810 187 837 209
819 194 827 210
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
202 1007 229 1029
211 1014 219 1030
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
196 1112 223 1134
205 1119 213 1135
1 K
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
377 1324 494 1346
387 1332 483 1348
12 JK Flip Flop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
377 591 396 615
382 595 390 611
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
383 791 402 815
388 795 396 811
1 K
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1064 336 1171 358
1073 344 1161 360
11 D Flip Flop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
372 357 503 379
381 365 493 381
14 D Flip Flop IC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
352 868 491 890
361 875 481 891
15 JK Flip Flop IC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
484 166 513 188
494 173 502 189
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
513 178 548 200
522 186 538 202
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1380 143 1409 165
1390 150 1398 166
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1387 227 1422 249
1396 235 1412 251
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
627 604 656 626
637 611 645 627
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
654 632 689 654
663 640 679 656
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
828 1038 857 1060
838 1045 846 1061
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
865 1060 900 1082
874 1068 890 1084
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
985 259 1010 281
993 266 1001 282
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
978 301 1013 323
987 308 1003 324
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1040 270 1063 292
1047 277 1055 293
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1167 145 1192 167
1175 153 1183 169
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1167 193 1192 215
1175 200 1183 216
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1223 162 1246 184
1230 169 1238 185
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1172 254 1207 276
1181 262 1197 278
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1172 290 1209 312
1182 298 1198 314
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1234 261 1269 283
1243 268 1259 284
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
351 1151 374 1173
358 1158 366 1174
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
351 1193 374 1215
358 1200 366 1216
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
395 1164 420 1186
403 1171 411 1187
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
474 1091 497 1113
481 1098 489 1114
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
473 1133 496 1155
480 1140 488 1156
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
516 1100 541 1122
524 1107 532 1123
1 3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
